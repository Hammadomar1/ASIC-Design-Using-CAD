module prbs_tb();

    timeunit 1ns;
    timeprecision 1ps;
    
    logic        data_in;
    logic        clk;
    logic        resetN;
    logic        load;
    logic        en;
    logic [1:15] seed = 15'b011011100010101;
    logic        ready_fec; // Ready from FEC
    logic        valid_in;  // Valid from testbench
    logic        data_out;
    logic        valid_out;
    logic        ready_randomizer; // Ready out from randomizer
    
    parameter CLK_PERIOD = 20;

    logic [95:0] data_in_sequence     = 96'hACBCD2114DAE1577C6DBF4C9;
    logic [95:0] data_out_expected    = 96'h558AC4A53A1724E163AC2BF9;
    logic [95:0] data_out_sequence;

    // ... [Clock generation and DUT instantiation remain the same]

    // Test sequence
    initial begin
        // Initialize signals
        resetN          = 0;
        load            = 0;
        en              = 0;
        valid_in        = 0;
        ready_fec       = 1;
        data_in         = 0;
        data_out_sequence = 0;

        // Reset sequence
        #(CLK_PERIOD);
        resetN = 1;
        #(CLK_PERIOD);

        // Load the seed
        load     = 1;
        en       = 0;
        valid_in = 0;
        #(CLK_PERIOD);
        load     = 0;

        // Enable PRBS operation
        en       = 1;
        valid_in = 1;
        #(CLK_PERIOD);

        // Wait for ready_randomizer
        wait (ready_randomizer == 1);

        // Send data sequence
        for (int i = 0; i < 96; i++) begin
            data_in = data_in_sequence[95 - i]; // Feeding from MSB to LSB
            #(CLK_PERIOD);
            data_out_sequence[95 - i] = data_out;
        end

        // Compare output with expected data
        if (data_out_sequence == data_out_expected) begin
            $display("Test passed");
        end else begin
            $display("Test failed");
            $display("Expected: %h", data_out_expected);
            $display("Got     : %h", data_out_sequence);
        end

        $stop();
    end
endmodule